-- Code your design here
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

-- Memória ROM 
-- Memória de instruções

entity mem_rom is
	generic (n: integer := 8; size: natural := 32);
	port (
	clock : in std_logic;
	address: in std_logic_vector(n-1 downto 0);
	dataout: out std_logic_vector(size - 1 downto 0)
	);
end mem_rom;

architecture RTL of mem_rom is 
type mem_type is array(0 to 31) of STD_LOGIC_VECTOR (31 downto 0);
signal mem: mem_type;
-- inicializando memória rom em  "00000000000000000000000000000000"
signal data_mem: mem_type := (

 	"00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 1
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 10 
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",  
        "00000000000000000000000000000000", -- mem 20
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 30
        "00000000000000000000000000000000"
);

begin 

dataout <= data_mem(to_integer(unsigned(address))) when (to_integer(unsigned(address))<((2**n)-1)) else (others => '0');


end RTL;